module registers;

endmodule
