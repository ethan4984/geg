`ifndef ALU_SVH_
`define ALU_SVH_ 

`define ALU_OP_ADD 0
`define ALU_OP_SUB 1

`endif
