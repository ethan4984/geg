`ifndef REGS_SVH_
`define REGS_SVH_

`define RF_PC 32

`endif
